module collision (
    input logic clk,
    input logic reset,
    input logic [9:0] bird_y,
    input logic [9:0] pipe_x,
    input logic [9:0] pipe_y_top,
    input logic [9:0] pipe_y_bot,

    output logic collided
);


endmodule