module prng (
    input logic clk,
    input logic reset,
    output logic [9:0] prng_out
);
assign prng_out = 500;

endmodule