`include "prng.sv"
`include "collision.sv"
module game_controller #(
    parameter int SCREEN_WIDTH    = 640, // Screen width in pixels
    parameter int SCREEN_HEIGHT   = 480, // Screen height in pixels
    parameter int PIPE_WIDTH      = 50,  // Pipe width in pixels
    parameter int PIPE_GAP        = 100, // Vertical gap between pipes
    parameter int PIPE_X_POS      = 300, // Horizontal position of the left edge of the pipes
    parameter int PIPE_GAP_Y_POS  = 190, // Vertical position of the top edge of the gap (0 = top)
    parameter int BIRD_WIDTH      = 20,  // Bird width in pixels
    parameter int BIRD_HEIGHT     = 20,  // Bird height in pixels
    // Calculate coordinate widths based on screen dimensions
    parameter int CORDW           = $clog2(SCREEN_WIDTH),
    parameter int CORDH           = $clog2(SCREEN_HEIGHT),
  	parameter logic [9:0] BIRD_X          = 500
) (
    input logic clk,
    input logic reset,
    input logic start_button,
    input logic [9:0] bird_y,
    // input logic [9:0] pipe_x,
    // input logic [9:0] pipe_y,
  	output logic collision_out,
    output logic [9:0] pipe_x_internal,
    output logic [9:0] pipe_y_bot,
    output logic [9:0] pipe_y_top
);
localparam logic [1:0] STATE_IDLE = 2'b00;
localparam logic [1:0] STATE_PLAY = 2'b01;
localparam logic [1:0] STATE_GAME_OVER = 2'b10;

logic [1:0] state;
logic [1:0] next_state;

// Declare internal signals for pipe position
logic [9:0] pipe_x_internal;
logic [9:0] pipe_y_internal;

logic [9:0] pipe_height;
//logic collision_out;

assign pipe_y_top = pipe_y_internal - PIPE_GAP;
assign pipe_y_bot = pipe_y_internal + PIPE_GAP;

always_ff @(posedge clk or negedge reset) begin
    if (reset) begin
        state <= STATE_IDLE;
    end
    else begin
        state <= next_state;
    end
end

always_ff @(posedge clk or negedge reset) begin
    if (reset) begin
        pipe_x_internal <= SCREEN_WIDTH;
        pipe_y_internal <= pipe_height;
    end
    else begin
        if (state == STATE_PLAY) begin
             if (pipe_x_internal > PIPE_WIDTH) begin
                 pipe_x_internal <= pipe_x_internal - 1;
             end else begin
                 pipe_x_internal <= SCREEN_WIDTH;
                 pipe_y_internal <= pipe_height;
             end
        end
    end
end

always_comb begin
    case (state)
        STATE_IDLE: begin
            if (start_button) begin
                next_state = STATE_PLAY;
            end
            else begin
                next_state = STATE_IDLE;
            end
        end
        STATE_PLAY: begin
            if (collision_out) begin
                next_state = STATE_GAME_OVER;
            end
            else begin
                next_state = STATE_PLAY;
            end
        end
        STATE_GAME_OVER: begin
            if (reset) begin
                next_state = STATE_IDLE;
            end
            else begin
                next_state = STATE_GAME_OVER;
            end
        end
        default: next_state = STATE_IDLE;
    endcase
end

// TODO: PRNG for pipe height generation
prng pipe_heights(.clk(clk), .reset(reset), .prng_out(pipe_height));

// TOOD: Collision module
collision collision_module(
    .clk(clk),
    .reset(reset),
    .bird_x(BIRD_X),
    .bird_y(bird_y),
    .pipe_x(pipe_x_internal),
    .pipe_y(pipe_y_internal),
    .collision_out(collision_out)
);

endmodule